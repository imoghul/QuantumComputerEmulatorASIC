    Mac OS X            	   2   �                                           ATTR         �   ,                  �     com.apple.quarantine    �     com.dropbox.attrs              com.dropbox.internal q/0081;00000000;; 

���]	�      WsϷ��	