    Mac OS X            	   2  
     <                                      ATTR      <      <                       com.apple.lastuseddate#PS           com.apple.quarantine   "     com.dropbox.attrs              com.dropbox.internal �re    x��$    q/0081;00000000;; 

���]	�      Wwֿ��	